module trn_cu(TxD_busy,clk,rst,FIR_valid,ff2_Sel,ff2_load,TxD_start);
input TxD_busy,clk,rst,FIR_valid;
output reg ff2_Sel,ff2_load,TxD_start;

reg [1:0]ns,ps;

parameter [1:0] idle=2'b00,
load_res=2'b01,
get_lsb=2'b10,
get_msb=2'b11;
always@(posedge clk)begin
    if(rst)
        {ff2_Sel,ff2_load,TxD_start,ns,ps}<=0;
    else begin
        ps<=ns;
    end
end
always@(*) begin
    case(ps)
    idle:ns=(FIR_valid==1'b1)?load_res:idle;
    load_res:ns=get_lsb;
    get_lsb:ns=(TxD_busy==1'b0)?get_msb:get_lsb;
    get_msb:ns=(TxD_busy==1'b0)?idle:get_msb;
endcase
end
always@(posedge clk) begin
     {ff2_Sel,ff2_load,TxD_start}=0;
    case(ps)
    idle:{ff2_load}=1'b1;
    load_res:{ff2_Sel,TxD_start}=2'b11;
    get_lsb:{TxD_start}=1'b0;
    get_msb:{ff2_Sel,TxD_start}=2'b01;
    endcase
end
endmodule