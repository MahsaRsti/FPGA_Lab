module CoefMem #(parameter width=16,length=64,adrlength=6) (
  rst,
  adr,
  d_out
  );
  input rst;
  input  [adrlength-1:0]   adr;
  output [width-1:0]   d_out;
  
  reg [width-1:0] mem[0:length-1];
  always @(posedge rst) begin
    mem[0] = 16'b0000000001111001;
    mem[1] = 16'b0000000001100000;
    mem[2] = 16'b1111111111001010;
    mem[3] = 16'b1111111011001010;
    mem[4] = 16'b1111111000011101;
    mem[5] = 16'b1111111001110101;
    mem[6] = 16'b1111111110110001;
    mem[7] = 16'b0000000011001010;
    mem[8] = 16'b0000000010111100;
    mem[9] = 16'b1111111110011110;
    mem[10] = 16'b1111111010110000;
    mem[11] = 16'b1111111100011110;
    mem[12] = 16'b0000000010100011;
    mem[13] = 16'b0000000110100010;
    mem[14] = 16'b0000000011010101;
    mem[15] = 16'b1111111011011110;
    mem[16] = 16'b1111110111100011;
    mem[17] = 16'b1111111101000101;
    mem[18] = 16'b0000000111010100;
    mem[19] = 16'b0000001010110011;
    mem[20] = 16'b0000000001110100;
    mem[21] = 16'b1111110100011100;
    mem[22] = 16'b1111110010000010;
    mem[23] = 16'b0000000000100000;
    mem[24] = 16'b0000010010110000;
    mem[25] = 16'b0000010010111111;
    mem[26] = 16'b1111111010001101;
    mem[27] = 16'b1111011101101001;
    mem[28] = 16'b1111100001010101;
    mem[29] = 16'b0000010111111001;
    mem[30] = 16'b0001101100000001;
    mem[31] = 16'b0010101011001000;
    mem[32] = 16'b0010101011001000;
    mem[33] = 16'b0001101100000001;
    mem[34] = 16'b0000010111111001;
    mem[35] = 16'b1111100001010101;
    mem[36] = 16'b1111011101101001;
    mem[37] = 16'b1111111010001101;
    mem[38] = 16'b0000010010111111;
    mem[39] = 16'b0000010010110000;
    mem[40] = 16'b0000000000100000;
    mem[41] = 16'b1111110010000010;
    mem[42] = 16'b1111110100011100;
    mem[43] = 16'b0000000001110100;
    mem[44] = 16'b0000001010110011;
    mem[45] = 16'b0000000111010100;
    mem[46] = 16'b1111111101000101;
    mem[47] = 16'b1111110111100011;
    mem[48] = 16'b1111111011011110;
    mem[49] = 16'b0000000011010101;
    mem[50] = 16'b0000000110100010;
    mem[51] = 16'b0000000010100011;
    mem[52] = 16'b1111111100011110;
    mem[53] = 16'b1111111010110000;
    mem[54] = 16'b1111111110011110;
    mem[55] = 16'b0000000010111100;
    mem[56] = 16'b0000000011001010;
    mem[57] = 16'b1111111110110001;
    mem[58] = 16'b1111111001110101;
    mem[59] = 16'b1111111000011101;
    mem[60] = 16'b1111111011001010;
    mem[61] = 16'b1111111111001010;
    mem[62] = 16'b0000000001100000;
    mem[63] = 16'b0000000001111001;
  end

  assign d_out = mem[adr];
  
endmodule   
